module stopwatch (
    input logic clk, nrst, pb0, pb1,
    output logic [6:0] out0, out1, out2, out3
);





endmodule